`include "svunit_defines.svh"
`include "svunit_assert_macros.svh"

module xcom_unit_test;
import svunit_pkg::svunit_testcase;

  string name = "xcom_ut";
  svunit_testcase svunit_ut;

  localparam CLOCK_FREQUENCY = 250e6; //[Hz]
  localparam SYNC_PULSE_FREQ = 5e6; //[Hz]

  localparam NB                 = 32;

  logic          tb_clk         = 1'b0;
  logic          tb_rstn        = 1'b1;
  logic          tb_i_sync      = 1'b0;
  logic [ 4-1:0] tb_i_cfg_tick  = 4'b0000;
  logic          tb_i_req       = 1'b0;
  logic          tb_i_valid     = 1'b0;
  logic [ 8-1:0] tb_i_header    = 8'b0000_0000;
  logic [NB-1:0] tb_i_data      = 32'h00000000; 
  logic          tb_o_ready     ;
  logic          tb_o_data      ;
  logic          tb_o_clk       ;
  logic [2-1:0]  tb_o_dbg_state ; 

initial begin
  $dumpfile("xcom.vcd");
  $dumpvars();
end

clk_gen
#(
  .FREQ       ( CLOCK_FREQUENCY   )
)
u_clk_gen
(
  .i_enable   ( 1'b1              ),
  .o_clk      ( tb_clk            )
);

clocking cb @(posedge tb_clk);
  default input #1step output #2;
  output  tb_rstn          ;
  output  tb_i_sync        ;
  output  tb_i_cfg_tick    ;
  output  tb_i_req         ;
  output  tb_i_valid       ;
  output  tb_i_header      ;
  output  tb_i_data        ;

  input   tb_o_ready       ;
  input   tb_o_data        ;
  input   tb_o_clk         ;
  input   tb_o_dbg_state   ;
endclocking

initial begin
  tb_i_sync <= 1'b0;
  forever # (200) tb_i_sync <= ~tb_i_sync;  
end 



//===================================
// This is the UUT that we're
// running the Unit Tests on
//===================================

xcom#(
   .NCH          ( 2 ), 
   .SYNC         ( 1 ), 
   .DEBUG        ( 1 )
) u_xcom(
   .i_ps_clk           ( tb_clk  ),   
   .i_ps_rstn          ( tb_rstn ),   
   .i_core_clk         (),   
   .i_core_rstn        (),   
   .i_time_clk         (),   
   .i_time_rstn        (),   
   .i_core_en          (),   
   .i_core_op          (),   
   .i_core_data1       (),   
   .i_core_data2       (),   
   .o_core_ready       (),   
   .o_core_data1       (),   
   .o_core_data2       (),   
   .o_core_valid       (),   
   .o_core_flag        (),   
   .i_sync             (),   
   .o_proc_start       (),   
   .o_proc_stop        (),   
   .o_time_rst         (),   
   .o_time_update      (),   
   .o_time_update_data (),
   .o_core_start       (),   
   .o_core_stop        (),   
   .o_xcom_id          (),   
   .i_xcom_clk         (),   
   .i_xcom_data        (),   
   .o_xcom_clk         (),   
   .o_xcom_data        (),   
   .s_axi_awaddr       (),   
   .s_axi_awprot       (),   
   .s_axi_awvalid      (),   
   .s_axi_awready      (),   
   .s_axi_wdata        (),   
   .s_axi_wstrb        (),   
   .s_axi_wvalid       (),   
   .s_axi_wready       (),   
   .s_axi_bresp        (),   
   .s_axi_bvalid       (),   
   .s_axi_bready       (),   
   .s_axi_araddr       (),   
   .s_axi_arprot       (),                                                                                                                                                                                             
   .s_axi_arvalid      (),   
   .s_axi_arready      (),   
   .s_axi_rdata        (),
   .s_axi_rresp        (),
   .s_axi_rvalid       (),
   .s_axi_rready       ()
);

//===================================
// Build
//===================================

function void build();
  svunit_ut = new(name);
endfunction

//===================================
// Setup for running the Unit Tests
//===================================
task setup();
  svunit_ut.setup();
    cb.tb_i_cfg_tick <= 4'h2;//N clock cycles in 1/0. Invalid values here 0 and 1. Bit LSB is always 0
    cb.tb_i_req      <= 1'b0;   
    cb.tb_i_valid    <= 1'b0;   
    cb.tb_i_header   <= 8'h00;   
    cb.tb_i_data     <= '0;

    @(cb);
    cb.tb_rstn    <= 1'b0;
    repeat(2) @(cb);
    cb.tb_rstn    <= 1'b1;
    repeat(5) @(cb);

endtask

//===================================
// Here we deconstruct anything we 
// need after running the Unit Tests
//===================================
task teardown();
  svunit_ut.teardown();
endtask

//===================================
// All tests are defined between the
// SVUNIT_TESTS_BEGIN/END macros
//
// Each individual test must be
// defined between `SVTEST(_NAME_)
// `SVTEST_END
//
// i.e.
//   `SVTEST(mytest)
//     <test code>
//   `SVTEST_END
//===================================

`SVUNIT_TESTS_BEGIN
`include "tests.sv"
`SVUNIT_TESTS_END 

endmodule
